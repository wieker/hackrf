module top(
    output IOB_0A, input IOB_6A
);

    assign IOB_0A = IOB_6A;

endmodule
